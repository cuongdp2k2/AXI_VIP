`ifndef LIB_SV
`define LIB_SV

`include"agent_active.sv"
`include"agent_passive.sv"
`include"base_env.sv"
`include"coverage.sv"
`include"driver.sv"
`include"env.sv"
`include"interface.sv"
`include"monitor.sv"
`include"package.sv"
`include"scoreboard.sv"
`include"seq_item.sv"
`include"sequence.sv"
`include"sequencer.sv"
`include"top.sv"

`endif 