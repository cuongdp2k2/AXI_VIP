interface B_IF(input CLK , RESET);
    logic [1:0]  BRESP  ;
    logic        BVALID ;
    logic        BREADY ;
endinterface //B_IF