interface IF (input clk , reset);

endinterface 